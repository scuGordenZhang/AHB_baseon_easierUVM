// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: AHB_slave_config.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-08-11 on Mon Jan 22 15:51:47 2018
//=============================================================================
// Description: Configuration for agent AHB_slave
//=============================================================================

`ifndef AHB_SLAVE_CONFIG_SV
`define AHB_SLAVE_CONFIG_SV

// You can insert code here by setting agent_config_inc_before_class in file AHB_slave.tpl

class AHB_slave_config extends uvm_object;

  // Do not register config class with the factory

  virtual AHB_slave_if     vif;
                  
  uvm_active_passive_enum  is_active = UVM_ACTIVE;
  bit                      coverage_enable;       
  bit                      checks_enable;         

  // You can insert variables here by setting config_var in file AHB_slave.tpl

  // You can remove new by setting agent_config_generate_methods_inside_class = no in file AHB_slave.tpl

  extern function new(string name = "");

  // You can insert code here by setting agent_config_inc_inside_class in file AHB_slave.tpl

endclass : AHB_slave_config 


// You can remove new by setting agent_config_generate_methods_after_class = no in file AHB_slave.tpl

function AHB_slave_config::new(string name = "");
  super.new(name);
endfunction : new


// You can insert code here by setting agent_config_inc_after_class in file AHB_slave.tpl

`endif // AHB_SLAVE_CONFIG_SV

