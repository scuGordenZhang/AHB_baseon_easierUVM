package sequences_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;
  import AHB_master_agent_pkg::*;

  `include "reset_seq.sv"

  `include "AHB_master_seq_lib.sv"

  

endpackage : sequences_pkg
