// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: AHB_master_sequencer.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-08-11 on Mon Jan 22 15:51:47 2018
//=============================================================================
// Description: Sequencer for AHB_master
//=============================================================================

`ifndef AHB_MASTER_SEQUENCER_SV
`define AHB_MASTER_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(trans) AHB_master_sequencer_t;


`endif // AHB_MASTER_SEQUENCER_SV

